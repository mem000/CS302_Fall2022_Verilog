-------------------------------------------------------------------------------
--
-- Title       : Prob_3_39
-- Design      : CS302_Fall2022
-- Author      : Mahmoud Esmat
-- Company     : MEM
--
-------------------------------------------------------------------------------
--
-- File        : F:\Verilog_Projects\ActHDL_Designs\CS302_Fall2022\CS302_Fall2022\src\Prob_3_39.vhd
-- Generated   : Sat Nov  5 01:27:57 2022
-- From        : interface description file
-- By          : Itf2Vhdl ver. 1.22
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------

--{{ Section below this comment is automatically maintained
--   and may be overwritten
--{entity {Prob_3_39} architecture {Prob_3_39}}



entity Prob_3_39 is
end Prob_3_39;

--}} End of automatically maintained section

architecture Prob_3_39 of Prob_3_39 is
begin

	 -- enter your statements here --

end Prob_3_39;
